* inverter

.subckt inverter in out

.param pmL=65n pmW=215n pmOX=1.95n nmL=65n nmW=130n nmOX=1.85n  

M1 out in vdd vdd tp L=pmL W=pmW
*                    L=65n  W=215n 

+ AS=75.3f AD=75.3f PS=1.23u PD=1.23u

M2 out in vss vss tn L=nmL W=nmW
*                    L=65n  W=130n 

+ AS=75.3f AD=75.3f PS=1.12u PD=1.23u

* BSIM4 4.8.2 models
* put here your .model statements from the previous question
.model tp pmos level=54 version=4.8.2 TOXE=pmOX
*                                     TOXE=1.95n

.model tn nmos level=54 version=4.8.2 TOXE=nmOX
*                                     TOXE=1.85n

.ends inverter




